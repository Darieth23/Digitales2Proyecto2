`include "Mux2a1_dest.v"
`include "Demux1a2_dest.v"
module enrrutamiento(
    //entradas


    //salidas



    );